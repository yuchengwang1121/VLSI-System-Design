

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO top 
  PIN ROM_address[11] 
    ANTENNAPARTIALMETALAREA 0.3948 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6356 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 0.6265 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 9.1504 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.2336 LAYER metal3 ;
  END ROM_address[11]
  PIN ROM_address[10] 
    ANTENNAPARTIALMETALAREA 149.884 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 620.948 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 0.6265 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 6.72 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1648 LAYER metal3 ;
  END ROM_address[10]
  PIN ROM_address[9] 
    ANTENNAPARTIALMETALAREA 8.3292 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.394 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 0.6265 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 28.2464 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 117.346 LAYER metal3 ;
  END ROM_address[9]
  PIN ROM_address[8] 
    ANTENNADIFFAREA 0.6265 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 154.202 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 639.16 LAYER metal2 ;
  END ROM_address[8]
  PIN ROM_address[7] 
    ANTENNADIFFAREA 1.0633 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 155.814 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 645.842 LAYER metal2 ;
  END ROM_address[7]
  PIN ROM_address[6] 
    ANTENNADIFFAREA 0.6265 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 160.082 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 663.52 LAYER metal2 ;
  END ROM_address[6]
  PIN ROM_address[5] 
    ANTENNADIFFAREA 0.6265 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 159.74 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 662.105 LAYER metal2 ;
  END ROM_address[5]
  PIN ROM_address[4] 
    ANTENNADIFFAREA 1.0633 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 159.076 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 659.356 LAYER metal2 ;
  END ROM_address[4]
  PIN ROM_address[3] 
    ANTENNADIFFAREA 1.0633 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 161.258 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 668.392 LAYER metal2 ;
  END ROM_address[3]
  PIN ROM_address[2] 
    ANTENNADIFFAREA 1.0633 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 161.798 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 670.631 LAYER metal2 ;
  END ROM_address[2]
  PIN ROM_address[1] 
    ANTENNADIFFAREA 0.5684 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 10.4552 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.964 LAYER metal2 ;
  END ROM_address[1]
  PIN ROM_address[0] 
    ANTENNADIFFAREA 1.0633 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 163.005 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 675.63 LAYER metal2 ;
  END ROM_address[0]
  PIN ROM_out[31] 
    ANTENNAPARTIALMETALAREA 7.9408 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.8976 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 54.782 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 227.279 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 53.7488 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 222.998 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 LAYER metal5 ; 
    ANTENNAMAXAREACAR 31.6014 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 134.324 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.59837 LAYER via5 ;
  END ROM_out[31]
  PIN ROM_out[30] 
    ANTENNAPARTIALMETALAREA 71.792 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 297.749 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3618 LAYER metal2 ; 
    ANTENNAMAXAREACAR 200.177 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 825.406 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.216694 LAYER via2 ;
  END ROM_out[30]
  PIN ROM_out[29] 
    ANTENNAPARTIALMETALAREA 4.9616 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5552 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 20.0228 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.2764 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 5.0176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.9472 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 24.9632 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1692.86 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5647.68 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5418.38 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18085.5 LAYER metal6 ;
  END ROM_out[29]
  PIN ROM_out[28] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.3612 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8212 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1732.51 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5779.84 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5541.79 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18494.3 LAYER metal6 ;
  END ROM_out[28]
  PIN ROM_out[27] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.3164 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6356 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1738.46 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5799.68 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5560.24 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18555.3 LAYER metal6 ;
  END ROM_out[27]
  PIN ROM_out[26] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2716 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.45 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1724.45 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5752.96 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5647.53 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18954.2 LAYER metal6 ;
  END ROM_out[26]
  PIN ROM_out[25] 
    ANTENNAPARTIALMETALAREA 5.0652 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.9844 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 30.8504 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 128.134 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 5.0176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 2.5424 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8576 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1695.55 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5656.64 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5425.52 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18108.1 LAYER metal6 ;
  END ROM_out[25]
  PIN ROM_out[24] 
    ANTENNAPARTIALMETALAREA 3.0736 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6208 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 18.3512 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.3512 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 13.1432 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 54.7752 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1713.02 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5714.88 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5487.72 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18321.7 LAYER metal6 ;
  END ROM_out[24]
  PIN ROM_out[23] 
    ANTENNAPARTIALMETALAREA 4.9756 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.6132 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 15.2264 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.4056 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.6704 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.6736 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.2032 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.5952 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1701.5 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5676.48 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5442.3 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18162.3 LAYER metal6 ;
  END ROM_out[23]
  PIN ROM_out[22] 
    ANTENNAPARTIALMETALAREA 5.3528 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0632 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 14.532 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.5288 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 5.0176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 7.336 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7168 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1694.88 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5654.4 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5426.09 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18112.2 LAYER metal6 ;
  END ROM_out[22]
  PIN ROM_out[21] 
    ANTENNAPARTIALMETALAREA 2.3128 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.5816 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 4.6368 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5344 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.6856 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.308 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1723.1 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5748.48 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5576.64 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18663 LAYER metal6 ;
  END ROM_out[21]
  PIN ROM_out[20] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 2.0832 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9552 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1729.15 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5768.64 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5543.08 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18508.3 LAYER metal6 ;
  END ROM_out[20]
  PIN ROM_out[19] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1735.2 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5788.8 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5551.95 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18529.4 LAYER metal6 ;
  END ROM_out[19]
  PIN ROM_out[18] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.6888 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1784 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1724.45 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5752.96 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5533.01 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18480.8 LAYER metal6 ;
  END ROM_out[18]
  PIN ROM_out[17] 
    ANTENNAPARTIALMETALAREA 3.5504 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7088 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.3892 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9372 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 13.7704 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 57.3736 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1721.76 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5744 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5509.37 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18387.8 LAYER metal6 ;
  END ROM_out[17]
  PIN ROM_out[16] 
    ANTENNAPARTIALMETALAREA 8.2544 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.1968 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 9.3856 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.208 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.064 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7328 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.8984 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.1896 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1697.57 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5663.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5429.81 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18120.7 LAYER metal6 ;
  END ROM_out[16]
  PIN ROM_out[15] 
    ANTENNAPARTIALMETALAREA 2.4528 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1616 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.3108 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6124 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 20.9552 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 87.1392 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1716.38 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5726.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5513.99 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18421.8 LAYER metal6 ;
  END ROM_out[15]
  PIN ROM_out[14] 
    ANTENNAPARTIALMETALAREA 3.0764 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6324 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 15.9208 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.2824 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.7504 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4336 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1743.12 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5824.8 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5574.14 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18631.5 LAYER metal6 ;
  END ROM_out[14]
  PIN ROM_out[13] 
    ANTENNAPARTIALMETALAREA 2.7664 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4608 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 12.0372 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.1932 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1738.42 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5809.12 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5587.32 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18699.3 LAYER metal6 ;
  END ROM_out[13]
  PIN ROM_out[12] 
    ANTENNAPARTIALMETALAREA 0.7504 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 7.7616 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.48 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1725.12 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5755.2 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5534.3 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18484.4 LAYER metal6 ;
  END ROM_out[12]
  PIN ROM_out[11] 
    ANTENNAPARTIALMETALAREA 0.364 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.508 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 9.5312 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.8112 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.7248 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.4704 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1704.14 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5694.88 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5470.71 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18305.8 LAYER metal6 ;
  END ROM_out[11]
  PIN ROM_out[10] 
    ANTENNAPARTIALMETALAREA 2.7664 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4608 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 5.7568 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.1744 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2736 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1717.06 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5728.32 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5528.26 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18478.2 LAYER metal6 ;
  END ROM_out[10]
  PIN ROM_out[9] 
    ANTENNAPARTIALMETALAREA 401.912 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1665.71 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 22.5008 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 93.5424 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 86.795 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 356.659 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[9]
  PIN ROM_out[8] 
    ANTENNAPARTIALMETALAREA 403.25 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1670.93 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.94317 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 25.8442 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[8]
  PIN ROM_out[7] 
    ANTENNAPARTIALMETALAREA 4.326 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.2212 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 18.5383 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 75.9553 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[7]
  PIN ROM_out[6] 
    ANTENNAPARTIALMETALAREA 141.252 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 585.51 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 18.4936 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 74.7331 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END ROM_out[6]
  PIN ROM_out[5] 
    ANTENNAPARTIALMETALAREA 141.246 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 585.487 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 24.5192 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 99.696 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END ROM_out[5]
  PIN ROM_out[4] 
    ANTENNAPARTIALMETALAREA 149.47 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 619.556 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.4216 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.5 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal5 ; 
    ANTENNAMAXAREACAR 33.03 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 137.029 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.00128 LAYER via5 ;
  END ROM_out[4]
  PIN ROM_out[3] 
    ANTENNAPARTIALMETALAREA 3.7324 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.762 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 16.9649 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 69.4368 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[3]
  PIN ROM_out[2] 
    ANTENNAPARTIALMETALAREA 176.54 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 731.705 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 18.9406 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 78.659 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END ROM_out[2]
  PIN ROM_out[1] 
    ANTENNAPARTIALMETALAREA 185.979 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 770.808 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 15.2931 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 63.5479 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END ROM_out[1]
  PIN ROM_out[0] 
    ANTENNAPARTIALMETALAREA 193.334 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 801.282 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.2896 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.096 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal5 ; 
    ANTENNAMAXAREACAR 237.451 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 981.844 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.00128 LAYER via5 ;
  END ROM_out[0]
  PIN DRAM_WEn[3] 
    ANTENNAPARTIALMETALAREA 204.814 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 848.517 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 5.20755 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 198.576 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 822.997 LAYER metal4 ;
  END DRAM_WEn[3]
  PIN DRAM_WEn[2] 
    ANTENNAPARTIALMETALAREA 205.713 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 852.24 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 5.20755 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 180.93 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 749.894 LAYER metal4 ;
  END DRAM_WEn[2]
  PIN DRAM_WEn[1] 
    ANTENNAPARTIALMETALAREA 206.175 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 854.154 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 5.20755 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 155.742 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 645.54 LAYER metal4 ;
  END DRAM_WEn[1]
  PIN DRAM_WEn[0] 
    ANTENNAPARTIALMETALAREA 115.29 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 477.63 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 4.8649 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 61.936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 256.917 LAYER metal4 ;
  END DRAM_WEn[0]
  PIN DRAM_A[10] 
    ANTENNAPARTIALMETALAREA 94.444 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 391.268 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 61.8856 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 256.708 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.28045 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 119.252 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 494.369 LAYER metal5 ;
  END DRAM_A[10]
  PIN DRAM_A[9] 
    ANTENNAPARTIALMETALAREA 144.872 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 600.184 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 35.14 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 145.905 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 66.2704 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 274.874 LAYER metal5 ;
  END DRAM_A[9]
  PIN DRAM_A[8] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.74 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.1616 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.28 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 211.882 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 878.12 LAYER metal5 ;
  END DRAM_A[8]
  PIN DRAM_A[7] 
    ANTENNAPARTIALMETALAREA 0.4872 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0184 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.0432 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0752 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 213.758 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 885.892 LAYER metal5 ;
  END DRAM_A[7]
  PIN DRAM_A[6] 
    ANTENNAPARTIALMETALAREA 0.4424 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8328 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.2208 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3824 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 213.097 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 883.154 LAYER metal5 ;
  END DRAM_A[6]
  PIN DRAM_A[5] 
    ANTENNAPARTIALMETALAREA 2.5956 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7532 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 19.5832 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 81.4552 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 211.327 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 875.823 LAYER metal5 ;
  END DRAM_A[5]
  PIN DRAM_A[4] 
    ANTENNAPARTIALMETALAREA 3.7268 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.4396 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 38.2256 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 158.688 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 208.947 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 865.963 LAYER metal5 ;
  END DRAM_A[4]
  PIN DRAM_A[3] 
    ANTENNAPARTIALMETALAREA 3.3124 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7228 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 59.7408 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 247.822 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 210.162 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 870.998 LAYER metal5 ;
  END DRAM_A[3]
  PIN DRAM_A[2] 
    ANTENNAPARTIALMETALAREA 1.1228 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6516 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 72.7216 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 301.6 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 213.097 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 883.154 LAYER metal5 ;
  END DRAM_A[2]
  PIN DRAM_A[1] 
    ANTENNAPARTIALMETALAREA 2.814 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.658 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 87.0072 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 360.783 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 209.591 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 868.631 LAYER metal5 ;
  END DRAM_A[1]
  PIN DRAM_A[0] 
    ANTENNAPARTIALMETALAREA 0.3528 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 109.726 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 454.906 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 204.938 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 849.352 LAYER metal5 ;
  END DRAM_A[0]
  PIN DRAM_D[31] 
    ANTENNAPARTIALMETALAREA 2.492 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.324 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 3.416 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4768 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 200.738 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 831.952 LAYER metal5 ;
  END DRAM_D[31]
  PIN DRAM_D[30] 
    ANTENNAPARTIALMETALAREA 2.6012 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7764 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 6.5856 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.608 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 90.7088 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 376.118 LAYER metal5 ;
  END DRAM_D[30]
  PIN DRAM_D[29] 
    ANTENNAPARTIALMETALAREA 3.388 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.036 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 50.1592 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 208.127 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 54.1128 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 224.506 LAYER metal5 ;
  END DRAM_D[29]
  PIN DRAM_D[28] 
    ANTENNAPARTIALMETALAREA 3.4636 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3492 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.7888 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 141.193 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 585.266 LAYER metal5 ;
  END DRAM_D[28]
  PIN DRAM_D[27] 
    ANTENNAPARTIALMETALAREA 2.2008 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1176 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 93.016 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 385.677 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 54.6168 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 226.594 LAYER metal5 ;
  END DRAM_D[27]
  PIN DRAM_D[26] 
    ANTENNAPARTIALMETALAREA 2.8308 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7276 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 115.926 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 480.588 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 53.9392 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 223.787 LAYER metal5 ;
  END DRAM_D[26]
  PIN DRAM_D[25] 
    ANTENNAPARTIALMETALAREA 3.808 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.776 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 132.216 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 548.077 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 52.724 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 218.753 LAYER metal5 ;
  END DRAM_D[25]
  PIN DRAM_D[24] 
    ANTENNAPARTIALMETALAREA 3.5532 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7204 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 101.102 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 419.178 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 207.749 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 860.998 LAYER metal5 ;
  END DRAM_D[24]
  PIN DRAM_D[23] 
    ANTENNAPARTIALMETALAREA 1.5624 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4728 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 123.525 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 512.07 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 209.905 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 869.93 LAYER metal5 ;
  END DRAM_D[23]
  PIN DRAM_D[22] 
    ANTENNAPARTIALMETALAREA 1.8452 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6444 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 201.365 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 834.55 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 197.669 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 819.238 LAYER metal5 ;
  END DRAM_D[22]
  PIN DRAM_D[21] 
    ANTENNAPARTIALMETALAREA 1.0528 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 161.941 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 671.222 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 212.733 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 881.646 LAYER metal5 ;
  END DRAM_D[21]
  PIN DRAM_D[20] 
    ANTENNAPARTIALMETALAREA 2.4108 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9876 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 198.632 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 823.229 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 205.962 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 853.598 LAYER metal5 ;
  END DRAM_D[20]
  PIN DRAM_D[19] 
    ANTENNAPARTIALMETALAREA 1.428 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.916 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 266.75 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1105.43 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 199.248 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 825.781 LAYER metal5 ;
  END DRAM_D[19]
  PIN DRAM_D[18] 
    ANTENNAPARTIALMETALAREA 0.392 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.624 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 282.083 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1168.96 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.4202 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 201.846 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 836.546 LAYER metal5 ;
  END DRAM_D[18]
  PIN DRAM_D[17] 
    ANTENNAPARTIALMETALAREA 3.2256 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3632 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 232.378 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 963.032 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.4202 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 196.448 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 814.181 LAYER metal5 ;
  END DRAM_D[17]
  PIN DRAM_D[16] 
    ANTENNAPARTIALMETALAREA 0.728 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3408 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 61.6224 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 255.618 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.6902 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 201.09 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 833.414 LAYER metal5 ;
  END DRAM_D[16]
  PIN DRAM_D[15] 
    ANTENNAPARTIALMETALAREA 7 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 29 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 127.198 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 527.29 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 391.714 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1623.14 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 2.94815 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 7.9352 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1992 LAYER metal5 ;
  END DRAM_D[15]
  PIN DRAM_D[14] 
    ANTENNAPARTIALMETALAREA 7.9408 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.8976 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 43.8228 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 181.876 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 387.733 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1606.65 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.6902 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 73.2088 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 303.618 LAYER metal5 ;
  END DRAM_D[14]
  PIN DRAM_D[13] 
    ANTENNAPARTIALMETALAREA 7.954 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.8396 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 88.7992 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 368.207 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.6902 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 379.596 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1572.94 LAYER metal4 ;
  END DRAM_D[13]
  PIN DRAM_D[12] 
    ANTENNAPARTIALMETALAREA 341.536 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1414.93 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 44.044 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 182.793 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 55.0872 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 228.543 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.6902 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 33.2808 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 138.202 LAYER metal5 ;
  END DRAM_D[12]
  PIN DRAM_D[11] 
    ANTENNAPARTIALMETALAREA 392.308 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1625.6 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.6902 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 14.2912 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.5312 LAYER metal3 ;
  END DRAM_D[11]
  PIN DRAM_D[10] 
    ANTENNAPARTIALMETALAREA 295.042 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1222.32 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 21.8232 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 90.7352 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.6902 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 105.42 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 437.065 LAYER metal4 ;
  END DRAM_D[10]
  PIN DRAM_D[9] 
    ANTENNAPARTIALMETALAREA 347.474 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1439.54 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 13.1432 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.7752 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.6902 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 45.2816 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 187.92 LAYER metal4 ;
  END DRAM_D[9]
  PIN DRAM_D[8] 
    ANTENNAPARTIALMETALAREA 375.382 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1555.48 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 8.092 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.8488 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.6902 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 25.1552 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 104.539 LAYER metal4 ;
  END DRAM_D[8]
  PIN DRAM_D[7] 
    ANTENNAPARTIALMETALAREA 7.3884 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.4964 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 28.5936 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 118.784 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.6902 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 405.451 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1680.05 LAYER metal4 ;
  END DRAM_D[7]
  PIN DRAM_D[6] 
    ANTENNAPARTIALMETALAREA 7.7196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.9812 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 18.5248 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.0704 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.5386 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 387.262 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1604.7 LAYER metal4 ;
  END DRAM_D[6]
  PIN DRAM_D[5] 
    ANTENNADIFFAREA 1.6902 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 395.464 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1639 LAYER metal2 ;
  END DRAM_D[5]
  PIN DRAM_D[4] 
    ANTENNADIFFAREA 1.6902 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 394.565 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1634.95 LAYER metal2 ;
  END DRAM_D[4]
  PIN DRAM_D[3] 
    ANTENNAPARTIALMETALAREA 394.834 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1635.74 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.5386 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 13.9944 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.3016 LAYER metal3 ;
  END DRAM_D[3]
  PIN DRAM_D[2] 
    ANTENNAPARTIALMETALAREA 390.608 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1618.23 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.5386 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 35.5208 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 147.482 LAYER metal3 ;
  END DRAM_D[2]
  PIN DRAM_D[1] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 390.113 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1616.83 LAYER metal2 ;
  END DRAM_D[1]
  PIN DRAM_D[0] 
    ANTENNAPARTIALMETALAREA 391.174 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1620.58 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.5386 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 79.9456 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 331.528 LAYER metal3 ;
  END DRAM_D[0]
  PIN DRAM_Q[31] 
    ANTENNAPARTIALMETALAREA 7 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 29 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 10.9452 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.6692 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 395.416 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1638.48 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.2304 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6432 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal5 ; 
    ANTENNAMAXAREACAR 36.7079 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 140.042 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.22347 LAYER via5 ;
  END DRAM_Q[31]
  PIN DRAM_Q[30] 
    ANTENNAPARTIALMETALAREA 3.2416 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3168 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 32.9336 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 136.764 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1731.02 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5784.48 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5438.05 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18175.8 LAYER metal6 ;
  END DRAM_Q[30]
  PIN DRAM_Q[29] 
    ANTENNAPARTIALMETALAREA 2.5696 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5328 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 35.0168 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 145.394 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1736.16 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5792 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5454.96 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18200.7 LAYER metal6 ;
  END DRAM_Q[29]
  PIN DRAM_Q[28] 
    ANTENNAPARTIALMETALAREA 3.3256 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.6648 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 16.0944 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.0016 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1726.46 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5759.68 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5412 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18060.7 LAYER metal6 ;
  END DRAM_Q[28]
  PIN DRAM_Q[27] 
    ANTENNAPARTIALMETALAREA 2.6536 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8808 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 5.6784 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8496 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1718.69 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5733.76 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5408.87 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18075.5 LAYER metal6 ;
  END DRAM_Q[27]
  PIN DRAM_Q[26] 
    ANTENNAPARTIALMETALAREA 3.5504 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7088 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 4.5724 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.2676 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1715.04 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5721.6 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5386.05 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 17968.3 LAYER metal6 ;
  END DRAM_Q[26]
  PIN DRAM_Q[25] 
    ANTENNAPARTIALMETALAREA 1.3552 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6144 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.1844 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2316 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 2.2064 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4656 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1720.42 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5739.52 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5405.71 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18036.7 LAYER metal6 ;
  END DRAM_Q[25]
  PIN DRAM_Q[24] 
    ANTENNAPARTIALMETALAREA 2.6928 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0432 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 20.7816 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 86.42 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1719.74 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5737.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5396.09 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18012.8 LAYER metal6 ;
  END DRAM_Q[24]
  PIN DRAM_Q[23] 
    ANTENNAPARTIALMETALAREA 2.4528 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1616 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 11.3372 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.2932 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.7504 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4336 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1717.06 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5728.32 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5389.45 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 17993.1 LAYER metal6 ;
  END DRAM_Q[23]
  PIN DRAM_Q[22] 
    ANTENNAPARTIALMETALAREA 2.6032 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.672 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 13.1432 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.7752 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1715.71 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5723.84 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5429.6 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18166.9 LAYER metal6 ;
  END DRAM_Q[22]
  PIN DRAM_Q[21] 
    ANTENNAPARTIALMETALAREA 2.296 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.512 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 3.7828 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9964 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1719.74 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5737.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5407.2 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18044 LAYER metal6 ;
  END DRAM_Q[21]
  PIN DRAM_Q[20] 
    ANTENNAPARTIALMETALAREA 2.6096 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8112 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.6748 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1204 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.8176 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.712 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1713.7 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5717.12 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5375.81 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 17943.6 LAYER metal6 ;
  END DRAM_Q[20]
  PIN DRAM_Q[19] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.9348 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3404 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1739.23 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5802.24 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5460.34 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18230.8 LAYER metal6 ;
  END DRAM_Q[19]
  PIN DRAM_Q[18] 
    ANTENNAPARTIALMETALAREA 4.2356 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.4348 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 12.2752 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.1792 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1716.38 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5726.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5385.75 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 17963.9 LAYER metal6 ;
  END DRAM_Q[18]
  PIN DRAM_Q[17] 
    ANTENNAPARTIALMETALAREA 3.43 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.21 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 29.8088 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 123.818 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1720.03 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5738.24 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5404.39 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18046.5 LAYER metal6 ;
  END DRAM_Q[17]
  PIN DRAM_Q[16] 
    ANTENNAPARTIALMETALAREA 4.4708 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4092 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 44.2176 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 183.512 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.7504 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4336 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.6856 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.308 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1716.38 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5726.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5396.35 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18006.6 LAYER metal6 ;
  END DRAM_Q[16]
  PIN DRAM_Q[15] 
    ANTENNAPARTIALMETALAREA 2.9504 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1104 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 59.4944 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 246.802 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1733.04 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5791.2 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5444.92 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18196.9 LAYER metal6 ;
  END DRAM_Q[15]
  PIN DRAM_Q[14] 
    ANTENNAPARTIALMETALAREA 3.9388 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.2052 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 86.7496 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 359.716 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1731.7 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5786.72 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5439.9 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18194.1 LAYER metal6 ;
  END DRAM_Q[14]
  PIN DRAM_Q[13] 
    ANTENNAPARTIALMETALAREA 4.7536 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5808 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 113.764 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 471.633 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.064 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7328 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1733.47 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5783.04 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5436.35 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18143.9 LAYER metal6 ;
  END DRAM_Q[13]
  PIN DRAM_Q[12] 
    ANTENNAPARTIALMETALAREA 3.5468 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.5812 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 99.4224 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 412.218 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1735.06 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5797.92 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5447.1 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18217.4 LAYER metal6 ;
  END DRAM_Q[12]
  PIN DRAM_Q[11] 
    ANTENNAPARTIALMETALAREA 4.2868 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7596 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 70.952 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 294.269 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.7504 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4336 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1745.81 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5833.76 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5472.22 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18291.3 LAYER metal6 ;
  END DRAM_Q[11]
  PIN DRAM_Q[10] 
    ANTENNAPARTIALMETALAREA 3.1024 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.8528 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 223.272 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 925.309 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1719.74 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5737.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5401.29 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18018.7 LAYER metal6 ;
  END DRAM_Q[10]
  PIN DRAM_Q[9] 
    ANTENNAPARTIALMETALAREA 3.8948 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.1356 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 193.273 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 801.026 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1732.8 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5780.8 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5426.11 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18104.2 LAYER metal6 ;
  END DRAM_Q[9]
  PIN DRAM_Q[8] 
    ANTENNAPARTIALMETALAREA 2.6228 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7532 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 251.115 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1040.66 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1719.74 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5737.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5407.52 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18059.2 LAYER metal6 ;
  END DRAM_Q[8]
  PIN DRAM_Q[7] 
    ANTENNAPARTIALMETALAREA 7.296 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1136 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 357.515 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1481.78 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 3.416 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4768 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal4 ; 
    ANTENNAMAXAREACAR 82.9717 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 330.425 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.23598 LAYER via4 ;
  END DRAM_Q[7]
  PIN DRAM_Q[6] 
    ANTENNAPARTIALMETALAREA 400.512 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1659.26 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.632 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2288 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3204 LAYER metal4 ; 
    ANTENNAMAXAREACAR 35.2572 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 132.005 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.978777 LAYER via4 ;
  END DRAM_Q[6]
  PIN DRAM_Q[5] 
    ANTENNAPARTIALMETALAREA 3.1612 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0964 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 2.2064 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4656 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal5 ; 
    ANTENNAMAXAREACAR 61.5695 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 254.975 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.96032 LAYER via5 ;
  END DRAM_Q[5]
  PIN DRAM_Q[4] 
    ANTENNAPARTIALMETALAREA 23.9148 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 99.4004 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 LAYER metal3 ; 
    ANTENNAMAXAREACAR 132.031 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 542.656 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.799185 LAYER via3 ;
  END DRAM_Q[4]
  PIN DRAM_Q[3] 
    ANTENNAPARTIALMETALAREA 0.4088 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6936 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 353.08 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1463.08 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal5 ; 
    ANTENNAMAXAREACAR 42.1813 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 164.269 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.23318 LAYER via5 ;
  END DRAM_Q[3]
  PIN DRAM_Q[2] 
    ANTENNAPARTIALMETALAREA 10.2788 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.2332 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 2.9008 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3424 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 LAYER metal5 ; 
    ANTENNAMAXAREACAR 28.527 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 116.946 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.59837 LAYER via5 ;
  END DRAM_Q[2]
  PIN DRAM_Q[1] 
    ANTENNAPARTIALMETALAREA 338.097 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1401.01 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.0432 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0752 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal4 ; 
    ANTENNAMAXAREACAR 52.9468 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 206.854 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.71424 LAYER via4 ;
  END DRAM_Q[1]
  PIN DRAM_Q[0] 
    ANTENNAPARTIALMETALAREA 3.0772 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0732 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal4 ; 
    ANTENNAMAXAREACAR 33.059 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 125.708 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.987103 LAYER via4 ;
  END DRAM_Q[0]
  PIN sensor_out[31] 
    ANTENNAPARTIALMETALAREA 6.4316 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.97 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.0048 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6304 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 13.5051 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 54.0664 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END sensor_out[31]
  PIN sensor_out[30] 
    ANTENNAPARTIALMETALAREA 1.7192 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1224 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 205.531 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 851.811 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 12.1805 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 51.9179 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[30]
  PIN sensor_out[29] 
    ANTENNAPARTIALMETALAREA 2.4164 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0108 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 173.858 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 720.592 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.1968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.504 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 59.7563 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 246.985 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[29]
  PIN sensor_out[28] 
    ANTENNAPARTIALMETALAREA 1.5288 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3336 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 151.592 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 628.349 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 19.584 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal6 ; 
    ANTENNAMAXAREACAR 175.943 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 658.167 LAYER metal6 ;
  END sensor_out[28]
  PIN sensor_out[27] 
    ANTENNAPARTIALMETALAREA 2.9316 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1452 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.1872 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2176 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal5 ; 
    ANTENNAMAXAREACAR 30.4732 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 129.548 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.00128 LAYER via5 ;
  END sensor_out[27]
  PIN sensor_out[26] 
    ANTENNAPARTIALMETALAREA 184.758 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 765.751 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.9424 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6576 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 62.9028 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 251.818 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[26]
  PIN sensor_out[25] 
    ANTENNAPARTIALMETALAREA 182.014 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 754.383 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal4 ; 
    ANTENNAMAXAREACAR 4.86628 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 19.2894 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.561605 LAYER via4 ;
  END sensor_out[25]
  PIN sensor_out[24] 
    ANTENNAPARTIALMETALAREA 3.0492 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9572 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.5136 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.024 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 38.6149 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 149.146 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[24]
  PIN sensor_out[23] 
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal3 ; 
    ANTENNAMAXAREACAR 368.569 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 1516.1 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.989899 LAYER via3 ;
  END sensor_out[23]
  PIN sensor_out[22] 
    ANTENNAPARTIALMETALAREA 3.0492 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9572 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.8104 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2536 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 60.7109 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 242.737 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[22]
  PIN sensor_out[21] 
    ANTENNAPARTIALMETALAREA 179.427 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 743.664 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 21.9987 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 82.3586 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[21]
  PIN sensor_out[20] 
    ANTENNAPARTIALMETALAREA 179.284 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 742.748 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 27.4785 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 105.061 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[20]
  PIN sensor_out[19] 
    ANTENNAPARTIALMETALAREA 179.281 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 742.736 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 61.7008 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 246.838 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[19]
  PIN sensor_out[18] 
    ANTENNAPARTIALMETALAREA 179.41 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 743.595 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 18.0391 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 65.9545 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[18]
  PIN sensor_out[17] 
    ANTENNAPARTIALMETALAREA 2.912 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3888 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4544 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 40.4179 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 162.768 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[17]
  PIN sensor_out[16] 
    ANTENNAPARTIALMETALAREA 2.142 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1988 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal3 ; 
    ANTENNAMAXAREACAR 216.567 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 886.376 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.989899 LAYER via3 ;
  END sensor_out[16]
  PIN sensor_out[15] 
    ANTENNAPARTIALMETALAREA 170.4 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 706.266 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.8104 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2536 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 64.9886 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 260.46 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[15]
  PIN sensor_out[14] 
    ANTENNAPARTIALMETALAREA 3.206 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.6068 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 7.5208 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.4824 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 80.2967 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 325.929 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[14]
  PIN sensor_out[13] 
    ANTENNAPARTIALMETALAREA 179.892 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 745.59 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 21.9987 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 82.3586 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[13]
  PIN sensor_out[12] 
    ANTENNAPARTIALMETALAREA 179.6 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 744.384 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.1328 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.096 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 38.5442 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 152.955 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[12]
  PIN sensor_out[11] 
    ANTENNAPARTIALMETALAREA 182.171 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 755.032 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 56.822 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 226.626 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[11]
  PIN sensor_out[10] 
    ANTENNAPARTIALMETALAREA 179.743 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 744.975 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 23.0947 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 86.899 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[10]
  PIN sensor_out[9] 
    ANTENNAPARTIALMETALAREA 1.4924 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5076 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 167.759 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 695.327 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 45.226 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 184.737 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[9]
  PIN sensor_out[8] 
    ANTENNAPARTIALMETALAREA 2.2456 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3032 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 212.901 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 882.342 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal5 ; 
    ANTENNAMAXAREACAR 79.6967 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 329.326 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.00128 LAYER via5 ;
  END sensor_out[8]
  PIN sensor_out[7] 
    ANTENNAPARTIALMETALAREA 0.9996 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1412 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 218.232 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 904.429 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 17.568 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 63.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 67.6074 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 258.271 LAYER metal6 ;
  END sensor_out[7]
  PIN sensor_out[6] 
    ANTENNAPARTIALMETALAREA 2.9484 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.2148 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 240.654 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 997.322 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 20.9924 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 90.7507 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[6]
  PIN sensor_out[5] 
    ANTENNAPARTIALMETALAREA 1.3916 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7652 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 251.003 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1040.2 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 23.9876 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 100.833 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[5]
  PIN sensor_out[4] 
    ANTENNAPARTIALMETALAREA 2.6124 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8228 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 287.571 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1191.69 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 15.999 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 67.5912 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[4]
  PIN sensor_out[3] 
    ANTENNAPARTIALMETALAREA 1.9236 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9692 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 309.333 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1281.85 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 29.2999 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 122.309 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[3]
  PIN sensor_out[2] 
    ANTENNAPARTIALMETALAREA 4.8244 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3116 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.4752 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5792 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal4 ; 
    ANTENNAMAXAREACAR 15.1872 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 60.9799 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.561605 LAYER via4 ;
  END sensor_out[2]
  PIN sensor_out[1] 
    ANTENNAPARTIALMETALAREA 1.2236 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0692 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 361.144 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1496.49 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal5 ; 
    ANTENNAMAXAREACAR 76.2995 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 315.252 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.00128 LAYER via5 ;
  END sensor_out[1]
  PIN sensor_out[0] 
    ANTENNAPARTIALMETALAREA 0.4144 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7168 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 376.006 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1558.07 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 16.0525 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 67.5148 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.2184 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9048 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 111.748 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 463.281 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 235.166 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 974.586 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6406 LAYER metal4 ; 
    ANTENNAMAXAREACAR 90.5378 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 370.284 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.0890707 LAYER via4 ;
  END clk
  PIN clk2 
    ANTENNAPARTIALMETALAREA 0.2576 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0672 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 218.198 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 904.614 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.3622 LAYER metal4 ; 
    ANTENNAMAXAREACAR 42.2313 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 170.11 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.0438626 LAYER via4 ;
  END clk2
  PIN rst 
    ANTENNAPARTIALMETALAREA 10.8836 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.414 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 LAYER metal2 ; 
    ANTENNAMAXAREACAR 58.5912 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 236.752 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.399592 LAYER via2 ;
  END rst
  PIN rst2 
    ANTENNAPARTIALMETALAREA 276.069 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1144.04 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 9.4304 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.3936 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 LAYER metal3 ; 
    ANTENNAMAXAREACAR 272.56 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 1124.09 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.799185 LAYER via3 ;
  END rst2
  PIN DRAM_valid 
    ANTENNAPARTIALMETALAREA 2.7244 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6116 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 5.1744 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7616 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.369 LAYER metal4 ; 
    ANTENNAMAXAREACAR 41.3366 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 166.784 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.637398 LAYER via4 ;
  END DRAM_valid
  PIN sensor_ready 
    ANTENNAPARTIALMETALAREA 0.8652 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5844 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 252.918 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1048.13 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 399.426 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1655.09 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 38.928 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 144.16 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6294 LAYER metal6 ; 
    ANTENNAMAXAREACAR 77.4514 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 282.984 LAYER metal6 ;
  END sensor_ready
  PIN ROM_enable 
    ANTENNADIFFAREA 1.0633 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 13.1152 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.3344 LAYER metal2 ;
  END ROM_enable
  PIN ROM_read 
    ANTENNADIFFAREA 1.0633 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 27.7088 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 115.118 LAYER metal2 ;
  END ROM_read
  PIN DRAM_CSn 
    ANTENNAPARTIALMETALAREA 216.465 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 896.784 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.0927 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 221.805 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 919.555 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0464 LAYER metal4 ; 
    ANTENNAMAXAREACAR 246.651 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 1018.82 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.24682 LAYER via4 ;
  END DRAM_CSn
  PIN DRAM_RASn 
    ANTENNAPARTIALMETALAREA 217.308 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 900.276 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.66835 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 101.73 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 421.776 LAYER metal4 ;
  END DRAM_RASn
  PIN DRAM_CASn 
    ANTENNAPARTIALMETALAREA 87.3124 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 361.723 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 76.4848 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 317.19 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.66835 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 126.314 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 523.624 LAYER metal5 ;
  END DRAM_CASn
  PIN sensor_en 
    ANTENNAPARTIALMETALAREA 3.5084 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.5348 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 455.157 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1885.97 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.329 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 405.395 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1679.82 LAYER metal5 ;
  END sensor_en
END top

END LIBRARY
